//-----------------------------------
// File Name    : image_processing.v
// Module Name  : ImageProcessing
// Project      : Box Sorter
// Author       : Valerian Ratu
// Date         : February 6, 2018
//-----------------------------------

module ImageDecoding(
    rst,
    clk,

    // Either FIFO inputs
    // or if using internal FIFO
    // use 

)